module datapath (
    ports
);
    
endmodule