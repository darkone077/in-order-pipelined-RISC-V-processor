module deex (
    ports
);
    
endmodule